module functionABCreduced(
  input logic a, b,
  output logic Y
  
);

	and(Y, a, b);

endmodule