module decimal7decoder(
input logic [3:0] A,
output [6:0] Y,
output [6:0] Z );

always_comb
  begin
    case(A)
4'b1000 : Y[6:0]  = 7'b0000000; //-8
4'b1001 : Y[6:0]  = 7'b1111000; //-7
4'b1010 : Y[6:0]  = 7'b0000010; //-6
4'b1011 : Y[6:0]  = 7'b0010010; //-5
4'b1100 : Y[6:0]  = 7'b0011001; //-4
4'b1101 : Y[6:0]  = 7'b0110000; //-3
4'b1110 : Y[6:0]  = 7'b0100100; //-2
4'b1111 : Y[6:0]  = 7'b1111001; //-1
4'b0000 : Y[6:0]  = 7'b1000000; //0
4'b0001 : Y[6:0]  = 7'b1111001; //1
4'b0010 : Y[6:0]  = 7'b0100100; //2
4'b0011 : Y[6:0]  = 7'b0110000; //3
4'b0100 : Y[6:0]  = 7'b0011001; //4
4'b0101 : Y[6:0]  = 7'b0010010; //5
4'b0110 : Y[6:0]  = 7'b0000010; //6
4'b0111 : Y[6:0]  = 7'b1111000; //7 
default : Y[6:0]=7'b1111111;
endcase
end

always_comb
begin
case(A)
4'b1000 : Z[6:0]  = 7'b0111111; //-8
4'b1001 : Z[6:0]  = 7'b0111111; //-7
4'b1010 : Z[6:0]  = 7'b0111111; //-6
4'b1011 : Z[6:0]  = 7'b0111111; //-5
4'b1100 : Z[6:0]  = 7'b0111111; //-4
4'b1101 : Z[6:0]  = 7'b0111111; //-3
4'b1110 : Z[6:0]  = 7'b0111111; //-2
4'b1111 : Z[6:0]  = 7'b0111111; //-1
default : Z[6:0]  = 7'b1111111;

endcase
end

               

endmodule

